library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package git_hash_pkg is
    constant GIT_HASH : std_logic_vector(159 downto 0) := x"b0a652e36ad3b74f600a62dcf8a8796ecede8400";
end package;
