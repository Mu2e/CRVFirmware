gtp_xcvr.vhd