-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.11
--  \   \         Application : Spartan-6 FPGA GTP Transceiver Wizard
--  /   /         Filename : mgt_usrclk_source.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module MGT_USRCLK_SOURCE (for use with GTP Transceivers)
-- Generated by Xilinx Spartan-6 FPGA GTP Transceiver Wizard
-- 
-- 
-- (c) Copyright 2009 - 2011 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************
entity MGT_USRCLK_SOURCE is
generic
(
    FREQUENCY_MODE     : string   := "LOW";
    DIVIDE_2           : boolean  := false;
    FEEDBACK           : string   := "1X"; 
    DIVIDE             : real     := 2.0
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    CLK2X_OUT               : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    FB_IN                   : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);

end MGT_USRCLK_SOURCE;

architecture RTL of MGT_USRCLK_SOURCE is
--*********************************Wire Declarations***************************

    signal not_connected_i          : std_logic_vector(15 downto 0);
    signal clkdv_i                  : std_logic;
    signal clk0_i                   : std_logic;
    signal clk2x_i                  : std_logic;
    signal tied_to_ground_i         : std_logic;
    signal tied_to_ground_vec_i     : std_logic_vector(63 downto 0);

begin

--*********************************** Main Body of Code ***********************


    --  Static signal Assigments    
    tied_to_ground_i                  <= '0';        
    tied_to_ground_vec_i(63 downto 0) <= (others => '0');

    -- Instantiate a DCM module to divide the reference clock.
    clock_divider_i : DCM_SP
    generic map
    (
        CLKDV_DIVIDE          =>          DIVIDE,
        DFS_FREQUENCY_MODE    =>          "LOW", 
        CLKIN_DIVIDE_BY_2     =>          DIVIDE_2,
        CLK_FEEDBACK          =>          FEEDBACK,
        DLL_FREQUENCY_MODE    =>          FREQUENCY_MODE
    )    
    port map
    (
        CLK0                =>          clk0_i,
        CLK180              =>          open,
        CLK270              =>          open,
        CLK2X               =>          clk2x_i,
        CLK2X180            =>          open,
        CLK90               =>          open,
        CLKDV               =>          clkdv_i,
        CLKFX               =>          open,
        CLKFX180            =>          open,
        PSDONE              =>          open,
        STATUS              =>          open,
        DSSEN               =>          tied_to_ground_i,
        PSCLK               =>          tied_to_ground_i,
        PSEN                =>          tied_to_ground_i,          
        PSINCDEC            =>          tied_to_ground_i,      
        LOCKED              =>          DCM_LOCKED_OUT,
        CLKFB               =>          FB_IN,
        CLKIN               =>          CLK_IN,
        RST                 =>          DCM_RESET_IN
    );


    dcm_1x_bufg_i : BUFG
    port map
    (
        I                   =>          clk0_i,
        O                   =>          DIV1_OUT
    );
    
    dcm_2x_bufg_i : BUFG
    port map
    (
        I                   =>          clk2x_i,
        O                   =>          CLK2X_OUT
    );

    dcm_div2_bufg_i : BUFG 
    port map
    (
        I                   =>          clkdv_i,
        O                   =>          DIV2_OUT
    );



end RTL;

